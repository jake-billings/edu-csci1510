** Profile: "4_1_Multiplexer_Test_Billings-Multiplexer_Test_Sim_Billings"  [ C:\Users\student\Desktop\CSCI Labs\Lab06a_Billings\Lab06a_Billings-PSpiceFiles\4_1_Multiplexer_Test_Billings\Multiplexer_Test_Sim_Billings.sim ] 

** Creating circuit file "Multiplexer_Test_Sim_Billings.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../lab06a_billings_multiplexer_test_stim.stl" 
* From [PSPICE NETLIST] section of C:\Users\student\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\4_1_Multiplexer_Test_Billings.net" 


.END
