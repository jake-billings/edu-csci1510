** Profile: "SCHEMATIC1-Simulation_Part2"  [ C:\Users\student\Desktop\CSCI Labs\Lab03_Billings\Lab03_Billings-PSpiceFiles\SCHEMATIC1\Simulation_Part2.sim ] 

** Creating circuit file "Simulation_Part2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\student\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 
.stmlib "C:\Users\student\Desktop\CSCI Labs\Lab03_Billings_old\wxyz_base_500hz_billings.stl" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
