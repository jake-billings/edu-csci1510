** Profile: "MYSTERY-MYSTERY_Sim"  [ C:\Users\student\Desktop\CSCI Labs\Lab05_Billings\lab05_billings-pspicefiles\mystery\mystery_sim.sim ] 

** Creating circuit file "MYSTERY_Sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../clear.stl" 
* From [PSPICE NETLIST] section of C:\Users\student\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\MYSTERY.net" 


.END
