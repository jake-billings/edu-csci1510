** Profile: "GATES_Billings-ANDinput"  [ c:\users\student\desktop\csci labs\lab1_billings\lab1_billings-pspicefiles\gates_billings\andinput.sim ] 

** Creating circuit file "ANDinput.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../input.stl" 
* From [PSPICE NETLIST] section of C:\Users\student\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\GATES_Billings.net" 


.END
